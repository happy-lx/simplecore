module core(
  input   clock,
  input   reset,
  output  io_result
);
  assign io_result = 1'h0;
endmodule
