module AND(
  input   io_a,
  input   io_b,
  output  io_c
);
  assign io_c = io_a & io_b; // @[AND.scala 14:8]
endmodule
