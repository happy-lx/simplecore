module Cpath(
  input         clock,
  input         reset,
  output [2:0]  io_c2d_cp_pc_sel,
  output [1:0]  io_c2d_cp_op1_sel,
  output [1:0]  io_c2d_cp_op2_sel,
  output [4:0]  io_c2d_cp_alu_sel,
  output        io_c2d_cp_reg_wen,
  output        io_c2d_cp_mem_en,
  output [2:0]  io_c2d_cp_mem_read_op,
  output [7:0]  io_c2d_cp_mem_write_mask,
  output        io_c2d_cp_mem_wen,
  output [2:0]  io_c2d_cp_alu_ext_sel,
  output [1:0]  io_c2d_cp_wb_sel,
  output [2:0]  io_c2d_cp_csr_op,
  output        io_c2d_hasexception,
  output        io_c2d_shouldstall,
  input  [31:0] io_d2c_instr,
  input         io_d2c_islt,
  input         io_d2c_isltu,
  input         io_d2c_iseq,
  input         io_d2c_isredir,
  output        io_imem_req_ready,
  input         io_imem_req_valid,
  input  [31:0] io_imem_req_bits_addr,
  input  [7:0]  io_imem_req_bits_mask,
  input  [2:0]  io_imem_req_bits_op,
  input  [63:0] io_imem_req_bits_wdata,
  input         io_imem_req_bits_memen,
  input         io_imem_req_bits_wen,
  input         io_imem_resp_ready,
  output        io_imem_resp_valid,
  output [63:0] io_imem_resp_bits_rdata,
  output        io_dmem_req_ready,
  input         io_dmem_req_valid,
  input  [31:0] io_dmem_req_bits_addr,
  input  [7:0]  io_dmem_req_bits_mask,
  input  [2:0]  io_dmem_req_bits_op,
  input  [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_req_bits_memen,
  input         io_dmem_req_bits_wen,
  input         io_dmem_resp_ready,
  output        io_dmem_resp_valid,
  output [63:0] io_dmem_resp_bits_rdata
);
  wire [31:0] _T = io_d2c_instr & 32'h7f; // @[Lookup.scala 31:38]
  wire  _T_1 = 32'h6f == _T; // @[Lookup.scala 31:38]
  wire [31:0] _T_2 = io_d2c_instr & 32'h707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 32'h2067 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 32'h3 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_7 = 32'h4003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_9 = 32'h3003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_11 = 32'h1003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 32'h5003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_15 = 32'h2003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_17 = 32'h6003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_19 = 32'h37 == _T; // @[Lookup.scala 31:38]
  wire  _T_21 = 32'h17 == _T; // @[Lookup.scala 31:38]
  wire [31:0] _T_22 = io_d2c_instr & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_23 = 32'h1033 == _T_22; // @[Lookup.scala 31:38]
  wire [31:0] _T_24 = io_d2c_instr & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_25 = 32'h101b == _T_24; // @[Lookup.scala 31:38]
  wire  _T_29 = 32'h103b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_31 = 32'h2033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_33 = 32'h2013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_35 = 32'h3013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_37 = 32'h3033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_39 = 32'h40005033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_41 = 32'h40005013 == _T_24; // @[Lookup.scala 31:38]
  wire  _T_43 = 32'h4000501b == _T_24; // @[Lookup.scala 31:38]
  wire  _T_45 = 32'h4000503b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_47 = 32'h5033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_49 = 32'h5013 == _T_24; // @[Lookup.scala 31:38]
  wire  _T_51 = 32'h501b == _T_24; // @[Lookup.scala 31:38]
  wire  _T_53 = 32'h503b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_55 = 32'h40000033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_57 = 32'h4000003b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_59 = 32'h4033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_61 = 32'h4013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_63 = 32'h33 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_65 = 32'h13 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_67 = 32'h1b == _T_2; // @[Lookup.scala 31:38]
  wire  _T_69 = 32'h3b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_71 = 32'h7033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_73 = 32'h7013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_75 = 32'h23 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_77 = 32'h3023 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_79 = 32'h1023 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_81 = 32'h2023 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_83 = 32'h63 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_85 = 32'h5063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_87 = 32'h7063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_89 = 32'h4063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_91 = 32'h6063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_93 = 32'h1063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_95 = 32'h3073 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_97 = 32'h7073 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_99 = 32'h2073 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_101 = 32'h6073 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_103 = 32'h1073 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_105 = 32'h5073 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_107 = 32'h105073 == io_d2c_instr; // @[Lookup.scala 31:38]
  wire  _T_109 = 32'h73 == io_d2c_instr; // @[Lookup.scala 31:38]
  wire  _T_111 = 32'h10500073 == io_d2c_instr; // @[Lookup.scala 31:38]
  wire  _T_113 = 32'h10200073 == io_d2c_instr; // @[Lookup.scala 31:38]
  wire  _T_115 = 32'h30200073 == io_d2c_instr; // @[Lookup.scala 31:38]
  wire [31:0] _T_116 = io_d2c_instr & 32'hf00fffff; // @[Lookup.scala 31:38]
  wire  _T_117 = 32'hf == _T_116; // @[Lookup.scala 31:38]
  wire  _T_119 = 32'h100f == io_d2c_instr; // @[Lookup.scala 31:38]
  wire  _T_121 = 32'h2000033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_123 = 32'h2001033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_125 = 32'h2002033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_127 = 32'h2003033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_129 = 32'h200003b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_131 = 32'h2006033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_133 = 32'h2007033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_135 = 32'h200703b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_137 = 32'h200603b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_139 = 32'h2004033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_141 = 32'h2005033 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_143 = 32'h200503b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_145 = 32'h200403b == _T_22; // @[Lookup.scala 31:38]
  wire  _T_147 = _T_143 | _T_145; // @[Lookup.scala 33:37]
  wire  _T_148 = _T_141 | _T_147; // @[Lookup.scala 33:37]
  wire  _T_149 = _T_139 | _T_148; // @[Lookup.scala 33:37]
  wire  _T_150 = _T_137 | _T_149; // @[Lookup.scala 33:37]
  wire  _T_151 = _T_135 | _T_150; // @[Lookup.scala 33:37]
  wire  _T_152 = _T_133 | _T_151; // @[Lookup.scala 33:37]
  wire  _T_153 = _T_131 | _T_152; // @[Lookup.scala 33:37]
  wire  _T_154 = _T_129 | _T_153; // @[Lookup.scala 33:37]
  wire  _T_155 = _T_127 | _T_154; // @[Lookup.scala 33:37]
  wire  _T_156 = _T_125 | _T_155; // @[Lookup.scala 33:37]
  wire  _T_157 = _T_123 | _T_156; // @[Lookup.scala 33:37]
  wire  _T_158 = _T_121 | _T_157; // @[Lookup.scala 33:37]
  wire  _T_159 = _T_119 | _T_158; // @[Lookup.scala 33:37]
  wire  _T_160 = _T_117 | _T_159; // @[Lookup.scala 33:37]
  wire  _T_161 = _T_115 | _T_160; // @[Lookup.scala 33:37]
  wire  _T_162 = _T_113 | _T_161; // @[Lookup.scala 33:37]
  wire  _T_163 = _T_111 | _T_162; // @[Lookup.scala 33:37]
  wire  _T_164 = _T_109 | _T_163; // @[Lookup.scala 33:37]
  wire  _T_165 = _T_107 | _T_164; // @[Lookup.scala 33:37]
  wire  _T_166 = _T_105 | _T_165; // @[Lookup.scala 33:37]
  wire  _T_167 = _T_103 | _T_166; // @[Lookup.scala 33:37]
  wire  _T_168 = _T_101 | _T_167; // @[Lookup.scala 33:37]
  wire  _T_169 = _T_99 | _T_168; // @[Lookup.scala 33:37]
  wire  _T_170 = _T_97 | _T_169; // @[Lookup.scala 33:37]
  wire  _T_171 = _T_95 | _T_170; // @[Lookup.scala 33:37]
  wire  _T_172 = _T_93 | _T_171; // @[Lookup.scala 33:37]
  wire  _T_173 = _T_91 | _T_172; // @[Lookup.scala 33:37]
  wire  _T_174 = _T_89 | _T_173; // @[Lookup.scala 33:37]
  wire  _T_175 = _T_87 | _T_174; // @[Lookup.scala 33:37]
  wire  _T_176 = _T_85 | _T_175; // @[Lookup.scala 33:37]
  wire  _T_177 = _T_83 | _T_176; // @[Lookup.scala 33:37]
  wire  _T_178 = _T_81 | _T_177; // @[Lookup.scala 33:37]
  wire  _T_179 = _T_79 | _T_178; // @[Lookup.scala 33:37]
  wire  _T_180 = _T_77 | _T_179; // @[Lookup.scala 33:37]
  wire  _T_181 = _T_75 | _T_180; // @[Lookup.scala 33:37]
  wire  _T_182 = _T_73 | _T_181; // @[Lookup.scala 33:37]
  wire  _T_183 = _T_71 | _T_182; // @[Lookup.scala 33:37]
  wire  _T_184 = _T_69 | _T_183; // @[Lookup.scala 33:37]
  wire  _T_185 = _T_67 | _T_184; // @[Lookup.scala 33:37]
  wire  _T_186 = _T_65 | _T_185; // @[Lookup.scala 33:37]
  wire  _T_187 = _T_63 | _T_186; // @[Lookup.scala 33:37]
  wire  _T_188 = _T_61 | _T_187; // @[Lookup.scala 33:37]
  wire  _T_189 = _T_59 | _T_188; // @[Lookup.scala 33:37]
  wire  _T_190 = _T_57 | _T_189; // @[Lookup.scala 33:37]
  wire  _T_191 = _T_55 | _T_190; // @[Lookup.scala 33:37]
  wire  _T_192 = _T_53 | _T_191; // @[Lookup.scala 33:37]
  wire  _T_193 = _T_51 | _T_192; // @[Lookup.scala 33:37]
  wire  _T_194 = _T_49 | _T_193; // @[Lookup.scala 33:37]
  wire  _T_195 = _T_47 | _T_194; // @[Lookup.scala 33:37]
  wire  _T_196 = _T_45 | _T_195; // @[Lookup.scala 33:37]
  wire  _T_197 = _T_43 | _T_196; // @[Lookup.scala 33:37]
  wire  _T_198 = _T_41 | _T_197; // @[Lookup.scala 33:37]
  wire  _T_199 = _T_39 | _T_198; // @[Lookup.scala 33:37]
  wire  _T_200 = _T_37 | _T_199; // @[Lookup.scala 33:37]
  wire  _T_201 = _T_35 | _T_200; // @[Lookup.scala 33:37]
  wire  _T_202 = _T_33 | _T_201; // @[Lookup.scala 33:37]
  wire  _T_203 = _T_31 | _T_202; // @[Lookup.scala 33:37]
  wire  _T_204 = _T_29 | _T_203; // @[Lookup.scala 33:37]
  wire  _T_205 = _T_25 | _T_204; // @[Lookup.scala 33:37]
  wire  _T_206 = _T_25 | _T_205; // @[Lookup.scala 33:37]
  wire  _T_207 = _T_23 | _T_206; // @[Lookup.scala 33:37]
  wire  _T_208 = _T_21 | _T_207; // @[Lookup.scala 33:37]
  wire  _T_209 = _T_19 | _T_208; // @[Lookup.scala 33:37]
  wire  _T_210 = _T_17 | _T_209; // @[Lookup.scala 33:37]
  wire  _T_211 = _T_15 | _T_210; // @[Lookup.scala 33:37]
  wire  _T_212 = _T_13 | _T_211; // @[Lookup.scala 33:37]
  wire  _T_213 = _T_11 | _T_212; // @[Lookup.scala 33:37]
  wire  _T_214 = _T_9 | _T_213; // @[Lookup.scala 33:37]
  wire  _T_215 = _T_7 | _T_214; // @[Lookup.scala 33:37]
  wire  _T_216 = _T_5 | _T_215; // @[Lookup.scala 33:37]
  wire  _T_217 = _T_3 | _T_216; // @[Lookup.scala 33:37]
  wire  cs_valid_inst = _T_1 | _T_217; // @[Lookup.scala 33:37]
  wire [3:0] _T_244 = _T_93 ? 4'h2 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_245 = _T_91 ? 4'h4 : _T_244; // @[Lookup.scala 33:37]
  wire [3:0] _T_246 = _T_89 ? 4'h3 : _T_245; // @[Lookup.scala 33:37]
  wire [3:0] _T_247 = _T_87 ? 4'h6 : _T_246; // @[Lookup.scala 33:37]
  wire [3:0] _T_248 = _T_85 ? 4'h5 : _T_247; // @[Lookup.scala 33:37]
  wire [3:0] _T_249 = _T_83 ? 4'h1 : _T_248; // @[Lookup.scala 33:37]
  wire [3:0] _T_250 = _T_81 ? 4'h0 : _T_249; // @[Lookup.scala 33:37]
  wire [3:0] _T_251 = _T_79 ? 4'h0 : _T_250; // @[Lookup.scala 33:37]
  wire [3:0] _T_252 = _T_77 ? 4'h0 : _T_251; // @[Lookup.scala 33:37]
  wire [3:0] _T_253 = _T_75 ? 4'h0 : _T_252; // @[Lookup.scala 33:37]
  wire [3:0] _T_254 = _T_73 ? 4'h0 : _T_253; // @[Lookup.scala 33:37]
  wire [3:0] _T_255 = _T_71 ? 4'h0 : _T_254; // @[Lookup.scala 33:37]
  wire [3:0] _T_256 = _T_69 ? 4'h0 : _T_255; // @[Lookup.scala 33:37]
  wire [3:0] _T_257 = _T_67 ? 4'h0 : _T_256; // @[Lookup.scala 33:37]
  wire [3:0] _T_258 = _T_65 ? 4'h0 : _T_257; // @[Lookup.scala 33:37]
  wire [3:0] _T_259 = _T_63 ? 4'h0 : _T_258; // @[Lookup.scala 33:37]
  wire [3:0] _T_260 = _T_61 ? 4'h0 : _T_259; // @[Lookup.scala 33:37]
  wire [3:0] _T_261 = _T_59 ? 4'h0 : _T_260; // @[Lookup.scala 33:37]
  wire [3:0] _T_262 = _T_57 ? 4'h0 : _T_261; // @[Lookup.scala 33:37]
  wire [3:0] _T_263 = _T_55 ? 4'h0 : _T_262; // @[Lookup.scala 33:37]
  wire [3:0] _T_264 = _T_53 ? 4'h0 : _T_263; // @[Lookup.scala 33:37]
  wire [3:0] _T_265 = _T_51 ? 4'h0 : _T_264; // @[Lookup.scala 33:37]
  wire [3:0] _T_266 = _T_49 ? 4'h0 : _T_265; // @[Lookup.scala 33:37]
  wire [3:0] _T_267 = _T_47 ? 4'h0 : _T_266; // @[Lookup.scala 33:37]
  wire [3:0] _T_268 = _T_45 ? 4'h0 : _T_267; // @[Lookup.scala 33:37]
  wire [3:0] _T_269 = _T_43 ? 4'h0 : _T_268; // @[Lookup.scala 33:37]
  wire [3:0] _T_270 = _T_41 ? 4'h0 : _T_269; // @[Lookup.scala 33:37]
  wire [3:0] _T_271 = _T_39 ? 4'h0 : _T_270; // @[Lookup.scala 33:37]
  wire [3:0] _T_272 = _T_37 ? 4'h0 : _T_271; // @[Lookup.scala 33:37]
  wire [3:0] _T_273 = _T_35 ? 4'h0 : _T_272; // @[Lookup.scala 33:37]
  wire [3:0] _T_274 = _T_33 ? 4'h0 : _T_273; // @[Lookup.scala 33:37]
  wire [3:0] _T_275 = _T_31 ? 4'h0 : _T_274; // @[Lookup.scala 33:37]
  wire [3:0] _T_276 = _T_29 ? 4'h0 : _T_275; // @[Lookup.scala 33:37]
  wire [3:0] _T_277 = _T_25 ? 4'h0 : _T_276; // @[Lookup.scala 33:37]
  wire [3:0] _T_278 = _T_25 ? 4'h0 : _T_277; // @[Lookup.scala 33:37]
  wire [3:0] _T_279 = _T_23 ? 4'h0 : _T_278; // @[Lookup.scala 33:37]
  wire [3:0] _T_280 = _T_21 ? 4'h0 : _T_279; // @[Lookup.scala 33:37]
  wire [3:0] _T_281 = _T_19 ? 4'h0 : _T_280; // @[Lookup.scala 33:37]
  wire [3:0] _T_282 = _T_17 ? 4'h0 : _T_281; // @[Lookup.scala 33:37]
  wire [3:0] _T_283 = _T_15 ? 4'h0 : _T_282; // @[Lookup.scala 33:37]
  wire [3:0] _T_284 = _T_13 ? 4'h0 : _T_283; // @[Lookup.scala 33:37]
  wire [3:0] _T_285 = _T_11 ? 4'h0 : _T_284; // @[Lookup.scala 33:37]
  wire [3:0] _T_286 = _T_9 ? 4'h0 : _T_285; // @[Lookup.scala 33:37]
  wire [3:0] _T_287 = _T_7 ? 4'h0 : _T_286; // @[Lookup.scala 33:37]
  wire [3:0] _T_288 = _T_5 ? 4'h0 : _T_287; // @[Lookup.scala 33:37]
  wire [3:0] _T_289 = _T_3 ? 4'h8 : _T_288; // @[Lookup.scala 33:37]
  wire [3:0] cs_branch = _T_1 ? 4'h7 : _T_289; // @[Lookup.scala 33:37]
  wire [1:0] _T_310 = _T_105 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_311 = _T_103 ? 2'h0 : _T_310; // @[Lookup.scala 33:37]
  wire [1:0] _T_312 = _T_101 ? 2'h1 : _T_311; // @[Lookup.scala 33:37]
  wire [1:0] _T_313 = _T_99 ? 2'h0 : _T_312; // @[Lookup.scala 33:37]
  wire [1:0] _T_314 = _T_97 ? 2'h1 : _T_313; // @[Lookup.scala 33:37]
  wire [1:0] _T_315 = _T_95 ? 2'h0 : _T_314; // @[Lookup.scala 33:37]
  wire [1:0] _T_316 = _T_93 ? 2'h0 : _T_315; // @[Lookup.scala 33:37]
  wire [1:0] _T_317 = _T_91 ? 2'h0 : _T_316; // @[Lookup.scala 33:37]
  wire [1:0] _T_318 = _T_89 ? 2'h0 : _T_317; // @[Lookup.scala 33:37]
  wire [1:0] _T_319 = _T_87 ? 2'h0 : _T_318; // @[Lookup.scala 33:37]
  wire [1:0] _T_320 = _T_85 ? 2'h0 : _T_319; // @[Lookup.scala 33:37]
  wire [1:0] _T_321 = _T_83 ? 2'h0 : _T_320; // @[Lookup.scala 33:37]
  wire [1:0] _T_322 = _T_81 ? 2'h0 : _T_321; // @[Lookup.scala 33:37]
  wire [1:0] _T_323 = _T_79 ? 2'h0 : _T_322; // @[Lookup.scala 33:37]
  wire [1:0] _T_324 = _T_77 ? 2'h0 : _T_323; // @[Lookup.scala 33:37]
  wire [1:0] _T_325 = _T_75 ? 2'h0 : _T_324; // @[Lookup.scala 33:37]
  wire [1:0] _T_326 = _T_73 ? 2'h0 : _T_325; // @[Lookup.scala 33:37]
  wire [1:0] _T_327 = _T_71 ? 2'h0 : _T_326; // @[Lookup.scala 33:37]
  wire [1:0] _T_328 = _T_69 ? 2'h0 : _T_327; // @[Lookup.scala 33:37]
  wire [1:0] _T_329 = _T_67 ? 2'h0 : _T_328; // @[Lookup.scala 33:37]
  wire [1:0] _T_330 = _T_65 ? 2'h0 : _T_329; // @[Lookup.scala 33:37]
  wire [1:0] _T_331 = _T_63 ? 2'h0 : _T_330; // @[Lookup.scala 33:37]
  wire [1:0] _T_332 = _T_61 ? 2'h0 : _T_331; // @[Lookup.scala 33:37]
  wire [1:0] _T_333 = _T_59 ? 2'h0 : _T_332; // @[Lookup.scala 33:37]
  wire [1:0] _T_334 = _T_57 ? 2'h0 : _T_333; // @[Lookup.scala 33:37]
  wire [1:0] _T_335 = _T_55 ? 2'h0 : _T_334; // @[Lookup.scala 33:37]
  wire [1:0] _T_336 = _T_53 ? 2'h0 : _T_335; // @[Lookup.scala 33:37]
  wire [1:0] _T_337 = _T_51 ? 2'h0 : _T_336; // @[Lookup.scala 33:37]
  wire [1:0] _T_338 = _T_49 ? 2'h0 : _T_337; // @[Lookup.scala 33:37]
  wire [1:0] _T_339 = _T_47 ? 2'h0 : _T_338; // @[Lookup.scala 33:37]
  wire [1:0] _T_340 = _T_45 ? 2'h0 : _T_339; // @[Lookup.scala 33:37]
  wire [1:0] _T_341 = _T_43 ? 2'h0 : _T_340; // @[Lookup.scala 33:37]
  wire [1:0] _T_342 = _T_41 ? 2'h0 : _T_341; // @[Lookup.scala 33:37]
  wire [1:0] _T_343 = _T_39 ? 2'h0 : _T_342; // @[Lookup.scala 33:37]
  wire [1:0] _T_344 = _T_37 ? 2'h0 : _T_343; // @[Lookup.scala 33:37]
  wire [1:0] _T_345 = _T_35 ? 2'h0 : _T_344; // @[Lookup.scala 33:37]
  wire [1:0] _T_346 = _T_33 ? 2'h0 : _T_345; // @[Lookup.scala 33:37]
  wire [1:0] _T_347 = _T_31 ? 2'h0 : _T_346; // @[Lookup.scala 33:37]
  wire [1:0] _T_348 = _T_29 ? 2'h0 : _T_347; // @[Lookup.scala 33:37]
  wire [1:0] _T_349 = _T_25 ? 2'h0 : _T_348; // @[Lookup.scala 33:37]
  wire [1:0] _T_350 = _T_25 ? 2'h0 : _T_349; // @[Lookup.scala 33:37]
  wire [1:0] _T_351 = _T_23 ? 2'h0 : _T_350; // @[Lookup.scala 33:37]
  wire [1:0] _T_352 = _T_21 ? 2'h2 : _T_351; // @[Lookup.scala 33:37]
  wire [1:0] _T_353 = _T_19 ? 2'h2 : _T_352; // @[Lookup.scala 33:37]
  wire [1:0] _T_354 = _T_17 ? 2'h0 : _T_353; // @[Lookup.scala 33:37]
  wire [1:0] _T_355 = _T_15 ? 2'h0 : _T_354; // @[Lookup.scala 33:37]
  wire [1:0] _T_356 = _T_13 ? 2'h0 : _T_355; // @[Lookup.scala 33:37]
  wire [1:0] _T_357 = _T_11 ? 2'h0 : _T_356; // @[Lookup.scala 33:37]
  wire [1:0] _T_358 = _T_9 ? 2'h0 : _T_357; // @[Lookup.scala 33:37]
  wire [1:0] _T_359 = _T_7 ? 2'h0 : _T_358; // @[Lookup.scala 33:37]
  wire [1:0] _T_360 = _T_5 ? 2'h0 : _T_359; // @[Lookup.scala 33:37]
  wire [1:0] _T_361 = _T_3 ? 2'h0 : _T_360; // @[Lookup.scala 33:37]
  wire [1:0] _T_394 = _T_81 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_395 = _T_79 ? 2'h3 : _T_394; // @[Lookup.scala 33:37]
  wire [1:0] _T_396 = _T_77 ? 2'h3 : _T_395; // @[Lookup.scala 33:37]
  wire [1:0] _T_397 = _T_75 ? 2'h3 : _T_396; // @[Lookup.scala 33:37]
  wire [1:0] _T_398 = _T_73 ? 2'h2 : _T_397; // @[Lookup.scala 33:37]
  wire [1:0] _T_399 = _T_71 ? 2'h0 : _T_398; // @[Lookup.scala 33:37]
  wire [1:0] _T_400 = _T_69 ? 2'h0 : _T_399; // @[Lookup.scala 33:37]
  wire [1:0] _T_401 = _T_67 ? 2'h2 : _T_400; // @[Lookup.scala 33:37]
  wire [1:0] _T_402 = _T_65 ? 2'h2 : _T_401; // @[Lookup.scala 33:37]
  wire [1:0] _T_403 = _T_63 ? 2'h0 : _T_402; // @[Lookup.scala 33:37]
  wire [1:0] _T_404 = _T_61 ? 2'h2 : _T_403; // @[Lookup.scala 33:37]
  wire [1:0] _T_405 = _T_59 ? 2'h0 : _T_404; // @[Lookup.scala 33:37]
  wire [1:0] _T_406 = _T_57 ? 2'h0 : _T_405; // @[Lookup.scala 33:37]
  wire [1:0] _T_407 = _T_55 ? 2'h0 : _T_406; // @[Lookup.scala 33:37]
  wire [1:0] _T_408 = _T_53 ? 2'h0 : _T_407; // @[Lookup.scala 33:37]
  wire [1:0] _T_409 = _T_51 ? 2'h2 : _T_408; // @[Lookup.scala 33:37]
  wire [1:0] _T_410 = _T_49 ? 2'h2 : _T_409; // @[Lookup.scala 33:37]
  wire [1:0] _T_411 = _T_47 ? 2'h0 : _T_410; // @[Lookup.scala 33:37]
  wire [1:0] _T_412 = _T_45 ? 2'h0 : _T_411; // @[Lookup.scala 33:37]
  wire [1:0] _T_413 = _T_43 ? 2'h2 : _T_412; // @[Lookup.scala 33:37]
  wire [1:0] _T_414 = _T_41 ? 2'h2 : _T_413; // @[Lookup.scala 33:37]
  wire [1:0] _T_415 = _T_39 ? 2'h0 : _T_414; // @[Lookup.scala 33:37]
  wire [1:0] _T_416 = _T_37 ? 2'h0 : _T_415; // @[Lookup.scala 33:37]
  wire [1:0] _T_417 = _T_35 ? 2'h2 : _T_416; // @[Lookup.scala 33:37]
  wire [1:0] _T_418 = _T_33 ? 2'h2 : _T_417; // @[Lookup.scala 33:37]
  wire [1:0] _T_419 = _T_31 ? 2'h0 : _T_418; // @[Lookup.scala 33:37]
  wire [1:0] _T_420 = _T_29 ? 2'h0 : _T_419; // @[Lookup.scala 33:37]
  wire [1:0] _T_421 = _T_25 ? 2'h2 : _T_420; // @[Lookup.scala 33:37]
  wire [1:0] _T_422 = _T_25 ? 2'h2 : _T_421; // @[Lookup.scala 33:37]
  wire [1:0] _T_423 = _T_23 ? 2'h0 : _T_422; // @[Lookup.scala 33:37]
  wire [1:0] _T_424 = _T_21 ? 2'h1 : _T_423; // @[Lookup.scala 33:37]
  wire [1:0] _T_425 = _T_19 ? 2'h0 : _T_424; // @[Lookup.scala 33:37]
  wire [1:0] _T_426 = _T_17 ? 2'h2 : _T_425; // @[Lookup.scala 33:37]
  wire [1:0] _T_427 = _T_15 ? 2'h2 : _T_426; // @[Lookup.scala 33:37]
  wire [1:0] _T_428 = _T_13 ? 2'h2 : _T_427; // @[Lookup.scala 33:37]
  wire [1:0] _T_429 = _T_11 ? 2'h2 : _T_428; // @[Lookup.scala 33:37]
  wire [1:0] _T_430 = _T_9 ? 2'h2 : _T_429; // @[Lookup.scala 33:37]
  wire [1:0] _T_431 = _T_7 ? 2'h2 : _T_430; // @[Lookup.scala 33:37]
  wire [1:0] _T_432 = _T_5 ? 2'h2 : _T_431; // @[Lookup.scala 33:37]
  wire [1:0] _T_433 = _T_3 ? 2'h0 : _T_432; // @[Lookup.scala 33:37]
  wire [4:0] _T_434 = _T_145 ? 5'h18 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_435 = _T_143 ? 5'h17 : _T_434; // @[Lookup.scala 33:37]
  wire [4:0] _T_436 = _T_141 ? 5'h16 : _T_435; // @[Lookup.scala 33:37]
  wire [4:0] _T_437 = _T_139 ? 5'h15 : _T_436; // @[Lookup.scala 33:37]
  wire [4:0] _T_438 = _T_137 ? 5'h14 : _T_437; // @[Lookup.scala 33:37]
  wire [4:0] _T_439 = _T_135 ? 5'h13 : _T_438; // @[Lookup.scala 33:37]
  wire [4:0] _T_440 = _T_133 ? 5'h12 : _T_439; // @[Lookup.scala 33:37]
  wire [4:0] _T_441 = _T_131 ? 5'h11 : _T_440; // @[Lookup.scala 33:37]
  wire [4:0] _T_442 = _T_129 ? 5'hd : _T_441; // @[Lookup.scala 33:37]
  wire [4:0] _T_443 = _T_127 ? 5'h10 : _T_442; // @[Lookup.scala 33:37]
  wire [4:0] _T_444 = _T_125 ? 5'hf : _T_443; // @[Lookup.scala 33:37]
  wire [4:0] _T_445 = _T_123 ? 5'he : _T_444; // @[Lookup.scala 33:37]
  wire [4:0] _T_446 = _T_121 ? 5'hd : _T_445; // @[Lookup.scala 33:37]
  wire [4:0] _T_447 = _T_119 ? 5'h0 : _T_446; // @[Lookup.scala 33:37]
  wire [4:0] _T_448 = _T_117 ? 5'h0 : _T_447; // @[Lookup.scala 33:37]
  wire [4:0] _T_449 = _T_115 ? 5'h0 : _T_448; // @[Lookup.scala 33:37]
  wire [4:0] _T_450 = _T_113 ? 5'h0 : _T_449; // @[Lookup.scala 33:37]
  wire [4:0] _T_451 = _T_111 ? 5'h0 : _T_450; // @[Lookup.scala 33:37]
  wire [4:0] _T_452 = _T_109 ? 5'h0 : _T_451; // @[Lookup.scala 33:37]
  wire [4:0] _T_453 = _T_107 ? 5'h0 : _T_452; // @[Lookup.scala 33:37]
  wire [4:0] _T_454 = _T_105 ? 5'hc : _T_453; // @[Lookup.scala 33:37]
  wire [4:0] _T_455 = _T_103 ? 5'hc : _T_454; // @[Lookup.scala 33:37]
  wire [4:0] _T_456 = _T_101 ? 5'hc : _T_455; // @[Lookup.scala 33:37]
  wire [4:0] _T_457 = _T_99 ? 5'hc : _T_456; // @[Lookup.scala 33:37]
  wire [4:0] _T_458 = _T_97 ? 5'hc : _T_457; // @[Lookup.scala 33:37]
  wire [4:0] _T_459 = _T_95 ? 5'hc : _T_458; // @[Lookup.scala 33:37]
  wire [4:0] _T_460 = _T_93 ? 5'h0 : _T_459; // @[Lookup.scala 33:37]
  wire [4:0] _T_461 = _T_91 ? 5'h0 : _T_460; // @[Lookup.scala 33:37]
  wire [4:0] _T_462 = _T_89 ? 5'h0 : _T_461; // @[Lookup.scala 33:37]
  wire [4:0] _T_463 = _T_87 ? 5'h0 : _T_462; // @[Lookup.scala 33:37]
  wire [4:0] _T_464 = _T_85 ? 5'h0 : _T_463; // @[Lookup.scala 33:37]
  wire [4:0] _T_465 = _T_83 ? 5'h0 : _T_464; // @[Lookup.scala 33:37]
  wire [4:0] _T_466 = _T_81 ? 5'h0 : _T_465; // @[Lookup.scala 33:37]
  wire [4:0] _T_467 = _T_79 ? 5'h0 : _T_466; // @[Lookup.scala 33:37]
  wire [4:0] _T_468 = _T_77 ? 5'h0 : _T_467; // @[Lookup.scala 33:37]
  wire [4:0] _T_469 = _T_75 ? 5'h0 : _T_468; // @[Lookup.scala 33:37]
  wire [4:0] _T_470 = _T_73 ? 5'h2 : _T_469; // @[Lookup.scala 33:37]
  wire [4:0] _T_471 = _T_71 ? 5'h2 : _T_470; // @[Lookup.scala 33:37]
  wire [4:0] _T_472 = _T_69 ? 5'h0 : _T_471; // @[Lookup.scala 33:37]
  wire [4:0] _T_473 = _T_67 ? 5'h0 : _T_472; // @[Lookup.scala 33:37]
  wire [4:0] _T_474 = _T_65 ? 5'h0 : _T_473; // @[Lookup.scala 33:37]
  wire [4:0] _T_475 = _T_63 ? 5'h0 : _T_474; // @[Lookup.scala 33:37]
  wire [4:0] _T_476 = _T_61 ? 5'h4 : _T_475; // @[Lookup.scala 33:37]
  wire [4:0] _T_477 = _T_59 ? 5'h4 : _T_476; // @[Lookup.scala 33:37]
  wire [4:0] _T_478 = _T_57 ? 5'h1 : _T_477; // @[Lookup.scala 33:37]
  wire [4:0] _T_479 = _T_55 ? 5'h1 : _T_478; // @[Lookup.scala 33:37]
  wire [4:0] _T_480 = _T_53 ? 5'hb : _T_479; // @[Lookup.scala 33:37]
  wire [4:0] _T_481 = _T_51 ? 5'hb : _T_480; // @[Lookup.scala 33:37]
  wire [4:0] _T_482 = _T_49 ? 5'ha : _T_481; // @[Lookup.scala 33:37]
  wire [4:0] _T_483 = _T_47 ? 5'ha : _T_482; // @[Lookup.scala 33:37]
  wire [4:0] _T_484 = _T_45 ? 5'h9 : _T_483; // @[Lookup.scala 33:37]
  wire [4:0] _T_485 = _T_43 ? 5'h9 : _T_484; // @[Lookup.scala 33:37]
  wire [4:0] _T_486 = _T_41 ? 5'h8 : _T_485; // @[Lookup.scala 33:37]
  wire [4:0] _T_487 = _T_39 ? 5'h8 : _T_486; // @[Lookup.scala 33:37]
  wire [4:0] _T_488 = _T_37 ? 5'h7 : _T_487; // @[Lookup.scala 33:37]
  wire [4:0] _T_489 = _T_35 ? 5'h7 : _T_488; // @[Lookup.scala 33:37]
  wire [4:0] _T_490 = _T_33 ? 5'h6 : _T_489; // @[Lookup.scala 33:37]
  wire [4:0] _T_491 = _T_31 ? 5'h6 : _T_490; // @[Lookup.scala 33:37]
  wire [4:0] _T_492 = _T_29 ? 5'h5 : _T_491; // @[Lookup.scala 33:37]
  wire [4:0] _T_493 = _T_25 ? 5'h5 : _T_492; // @[Lookup.scala 33:37]
  wire [4:0] _T_494 = _T_25 ? 5'h5 : _T_493; // @[Lookup.scala 33:37]
  wire [4:0] _T_495 = _T_23 ? 5'h5 : _T_494; // @[Lookup.scala 33:37]
  wire [4:0] _T_496 = _T_21 ? 5'h0 : _T_495; // @[Lookup.scala 33:37]
  wire [4:0] _T_497 = _T_19 ? 5'hc : _T_496; // @[Lookup.scala 33:37]
  wire [4:0] _T_498 = _T_17 ? 5'h0 : _T_497; // @[Lookup.scala 33:37]
  wire [4:0] _T_499 = _T_15 ? 5'h0 : _T_498; // @[Lookup.scala 33:37]
  wire [4:0] _T_500 = _T_13 ? 5'h0 : _T_499; // @[Lookup.scala 33:37]
  wire [4:0] _T_501 = _T_11 ? 5'h0 : _T_500; // @[Lookup.scala 33:37]
  wire [4:0] _T_502 = _T_9 ? 5'h0 : _T_501; // @[Lookup.scala 33:37]
  wire [4:0] _T_503 = _T_7 ? 5'h0 : _T_502; // @[Lookup.scala 33:37]
  wire [4:0] _T_504 = _T_5 ? 5'h0 : _T_503; // @[Lookup.scala 33:37]
  wire [4:0] _T_505 = _T_3 ? 5'h0 : _T_504; // @[Lookup.scala 33:37]
  wire  _T_519 = _T_119 ? 1'h0 : _T_158; // @[Lookup.scala 33:37]
  wire  _T_520 = _T_117 ? 1'h0 : _T_519; // @[Lookup.scala 33:37]
  wire  _T_521 = _T_115 ? 1'h0 : _T_520; // @[Lookup.scala 33:37]
  wire  _T_522 = _T_113 ? 1'h0 : _T_521; // @[Lookup.scala 33:37]
  wire  _T_523 = _T_111 ? 1'h0 : _T_522; // @[Lookup.scala 33:37]
  wire  _T_524 = _T_109 ? 1'h0 : _T_523; // @[Lookup.scala 33:37]
  wire  _T_525 = _T_107 ? 1'h0 : _T_524; // @[Lookup.scala 33:37]
  wire  _T_526 = _T_105 | _T_525; // @[Lookup.scala 33:37]
  wire  _T_527 = _T_103 | _T_526; // @[Lookup.scala 33:37]
  wire  _T_528 = _T_101 | _T_527; // @[Lookup.scala 33:37]
  wire  _T_529 = _T_99 | _T_528; // @[Lookup.scala 33:37]
  wire  _T_530 = _T_97 | _T_529; // @[Lookup.scala 33:37]
  wire  _T_531 = _T_95 | _T_530; // @[Lookup.scala 33:37]
  wire  _T_532 = _T_93 ? 1'h0 : _T_531; // @[Lookup.scala 33:37]
  wire  _T_533 = _T_91 ? 1'h0 : _T_532; // @[Lookup.scala 33:37]
  wire  _T_534 = _T_89 ? 1'h0 : _T_533; // @[Lookup.scala 33:37]
  wire  _T_535 = _T_87 ? 1'h0 : _T_534; // @[Lookup.scala 33:37]
  wire  _T_536 = _T_85 ? 1'h0 : _T_535; // @[Lookup.scala 33:37]
  wire  _T_537 = _T_83 ? 1'h0 : _T_536; // @[Lookup.scala 33:37]
  wire  _T_538 = _T_81 ? 1'h0 : _T_537; // @[Lookup.scala 33:37]
  wire  _T_539 = _T_79 ? 1'h0 : _T_538; // @[Lookup.scala 33:37]
  wire  _T_540 = _T_77 ? 1'h0 : _T_539; // @[Lookup.scala 33:37]
  wire  _T_541 = _T_75 ? 1'h0 : _T_540; // @[Lookup.scala 33:37]
  wire  _T_542 = _T_73 | _T_541; // @[Lookup.scala 33:37]
  wire  _T_543 = _T_71 | _T_542; // @[Lookup.scala 33:37]
  wire  _T_544 = _T_69 | _T_543; // @[Lookup.scala 33:37]
  wire  _T_545 = _T_67 | _T_544; // @[Lookup.scala 33:37]
  wire  _T_546 = _T_65 | _T_545; // @[Lookup.scala 33:37]
  wire  _T_547 = _T_63 | _T_546; // @[Lookup.scala 33:37]
  wire  _T_548 = _T_61 | _T_547; // @[Lookup.scala 33:37]
  wire  _T_549 = _T_59 | _T_548; // @[Lookup.scala 33:37]
  wire  _T_550 = _T_57 | _T_549; // @[Lookup.scala 33:37]
  wire  _T_551 = _T_55 | _T_550; // @[Lookup.scala 33:37]
  wire  _T_552 = _T_53 | _T_551; // @[Lookup.scala 33:37]
  wire  _T_553 = _T_51 | _T_552; // @[Lookup.scala 33:37]
  wire  _T_554 = _T_49 | _T_553; // @[Lookup.scala 33:37]
  wire  _T_555 = _T_47 | _T_554; // @[Lookup.scala 33:37]
  wire  _T_556 = _T_45 | _T_555; // @[Lookup.scala 33:37]
  wire  _T_557 = _T_43 | _T_556; // @[Lookup.scala 33:37]
  wire  _T_558 = _T_41 | _T_557; // @[Lookup.scala 33:37]
  wire  _T_559 = _T_39 | _T_558; // @[Lookup.scala 33:37]
  wire  _T_560 = _T_37 | _T_559; // @[Lookup.scala 33:37]
  wire  _T_561 = _T_35 | _T_560; // @[Lookup.scala 33:37]
  wire  _T_562 = _T_33 | _T_561; // @[Lookup.scala 33:37]
  wire  _T_563 = _T_31 | _T_562; // @[Lookup.scala 33:37]
  wire  _T_564 = _T_29 | _T_563; // @[Lookup.scala 33:37]
  wire  _T_565 = _T_25 | _T_564; // @[Lookup.scala 33:37]
  wire  _T_566 = _T_25 | _T_565; // @[Lookup.scala 33:37]
  wire  _T_567 = _T_23 | _T_566; // @[Lookup.scala 33:37]
  wire  _T_568 = _T_21 | _T_567; // @[Lookup.scala 33:37]
  wire  _T_569 = _T_19 | _T_568; // @[Lookup.scala 33:37]
  wire  _T_570 = _T_17 | _T_569; // @[Lookup.scala 33:37]
  wire  _T_571 = _T_15 | _T_570; // @[Lookup.scala 33:37]
  wire  _T_572 = _T_13 | _T_571; // @[Lookup.scala 33:37]
  wire  _T_573 = _T_11 | _T_572; // @[Lookup.scala 33:37]
  wire  _T_574 = _T_9 | _T_573; // @[Lookup.scala 33:37]
  wire  _T_575 = _T_7 | _T_574; // @[Lookup.scala 33:37]
  wire  _T_576 = _T_5 | _T_575; // @[Lookup.scala 33:37]
  wire  _T_577 = _T_3 ? 1'h0 : _T_576; // @[Lookup.scala 33:37]
  wire  _T_611 = _T_79 | _T_81; // @[Lookup.scala 33:37]
  wire  _T_612 = _T_77 | _T_611; // @[Lookup.scala 33:37]
  wire  _T_613 = _T_75 | _T_612; // @[Lookup.scala 33:37]
  wire  _T_614 = _T_73 ? 1'h0 : _T_613; // @[Lookup.scala 33:37]
  wire  _T_615 = _T_71 ? 1'h0 : _T_614; // @[Lookup.scala 33:37]
  wire  _T_616 = _T_69 ? 1'h0 : _T_615; // @[Lookup.scala 33:37]
  wire  _T_617 = _T_67 ? 1'h0 : _T_616; // @[Lookup.scala 33:37]
  wire  _T_618 = _T_65 ? 1'h0 : _T_617; // @[Lookup.scala 33:37]
  wire  _T_619 = _T_63 ? 1'h0 : _T_618; // @[Lookup.scala 33:37]
  wire  _T_620 = _T_61 ? 1'h0 : _T_619; // @[Lookup.scala 33:37]
  wire  _T_621 = _T_59 ? 1'h0 : _T_620; // @[Lookup.scala 33:37]
  wire  _T_622 = _T_57 ? 1'h0 : _T_621; // @[Lookup.scala 33:37]
  wire  _T_623 = _T_55 ? 1'h0 : _T_622; // @[Lookup.scala 33:37]
  wire  _T_624 = _T_53 ? 1'h0 : _T_623; // @[Lookup.scala 33:37]
  wire  _T_625 = _T_51 ? 1'h0 : _T_624; // @[Lookup.scala 33:37]
  wire  _T_626 = _T_49 ? 1'h0 : _T_625; // @[Lookup.scala 33:37]
  wire  _T_627 = _T_47 ? 1'h0 : _T_626; // @[Lookup.scala 33:37]
  wire  _T_628 = _T_45 ? 1'h0 : _T_627; // @[Lookup.scala 33:37]
  wire  _T_629 = _T_43 ? 1'h0 : _T_628; // @[Lookup.scala 33:37]
  wire  _T_630 = _T_41 ? 1'h0 : _T_629; // @[Lookup.scala 33:37]
  wire  _T_631 = _T_39 ? 1'h0 : _T_630; // @[Lookup.scala 33:37]
  wire  _T_632 = _T_37 ? 1'h0 : _T_631; // @[Lookup.scala 33:37]
  wire  _T_633 = _T_35 ? 1'h0 : _T_632; // @[Lookup.scala 33:37]
  wire  _T_634 = _T_33 ? 1'h0 : _T_633; // @[Lookup.scala 33:37]
  wire  _T_635 = _T_31 ? 1'h0 : _T_634; // @[Lookup.scala 33:37]
  wire  _T_636 = _T_29 ? 1'h0 : _T_635; // @[Lookup.scala 33:37]
  wire  _T_637 = _T_25 ? 1'h0 : _T_636; // @[Lookup.scala 33:37]
  wire  _T_638 = _T_25 ? 1'h0 : _T_637; // @[Lookup.scala 33:37]
  wire  _T_639 = _T_23 ? 1'h0 : _T_638; // @[Lookup.scala 33:37]
  wire  _T_640 = _T_21 ? 1'h0 : _T_639; // @[Lookup.scala 33:37]
  wire  _T_641 = _T_19 ? 1'h0 : _T_640; // @[Lookup.scala 33:37]
  wire  _T_642 = _T_17 | _T_641; // @[Lookup.scala 33:37]
  wire  _T_643 = _T_15 | _T_642; // @[Lookup.scala 33:37]
  wire  _T_644 = _T_13 | _T_643; // @[Lookup.scala 33:37]
  wire  _T_645 = _T_11 | _T_644; // @[Lookup.scala 33:37]
  wire  _T_646 = _T_9 | _T_645; // @[Lookup.scala 33:37]
  wire  _T_647 = _T_7 | _T_646; // @[Lookup.scala 33:37]
  wire  _T_648 = _T_5 | _T_647; // @[Lookup.scala 33:37]
  wire  _T_649 = _T_3 ? 1'h0 : _T_648; // @[Lookup.scala 33:37]
  wire [2:0] _T_714 = _T_17 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_715 = _T_15 ? 3'h4 : _T_714; // @[Lookup.scala 33:37]
  wire [2:0] _T_716 = _T_13 ? 3'h3 : _T_715; // @[Lookup.scala 33:37]
  wire [2:0] _T_717 = _T_11 ? 3'h2 : _T_716; // @[Lookup.scala 33:37]
  wire [2:0] _T_718 = _T_9 ? 3'h6 : _T_717; // @[Lookup.scala 33:37]
  wire [2:0] _T_719 = _T_7 ? 3'h1 : _T_718; // @[Lookup.scala 33:37]
  wire [2:0] _T_720 = _T_5 ? 3'h0 : _T_719; // @[Lookup.scala 33:37]
  wire [2:0] _T_721 = _T_3 ? 3'h0 : _T_720; // @[Lookup.scala 33:37]
  wire [7:0] _T_754 = _T_81 ? 8'h7 : 8'h1; // @[Lookup.scala 33:37]
  wire [7:0] _T_755 = _T_79 ? 8'h3 : _T_754; // @[Lookup.scala 33:37]
  wire [7:0] _T_756 = _T_77 ? 8'hf : _T_755; // @[Lookup.scala 33:37]
  wire [7:0] _T_757 = _T_75 ? 8'h1 : _T_756; // @[Lookup.scala 33:37]
  wire [7:0] _T_758 = _T_73 ? 8'h1 : _T_757; // @[Lookup.scala 33:37]
  wire [7:0] _T_759 = _T_71 ? 8'h1 : _T_758; // @[Lookup.scala 33:37]
  wire [7:0] _T_760 = _T_69 ? 8'h1 : _T_759; // @[Lookup.scala 33:37]
  wire [7:0] _T_761 = _T_67 ? 8'h1 : _T_760; // @[Lookup.scala 33:37]
  wire [7:0] _T_762 = _T_65 ? 8'h1 : _T_761; // @[Lookup.scala 33:37]
  wire [7:0] _T_763 = _T_63 ? 8'h1 : _T_762; // @[Lookup.scala 33:37]
  wire [7:0] _T_764 = _T_61 ? 8'h1 : _T_763; // @[Lookup.scala 33:37]
  wire [7:0] _T_765 = _T_59 ? 8'h1 : _T_764; // @[Lookup.scala 33:37]
  wire [7:0] _T_766 = _T_57 ? 8'h1 : _T_765; // @[Lookup.scala 33:37]
  wire [7:0] _T_767 = _T_55 ? 8'h1 : _T_766; // @[Lookup.scala 33:37]
  wire [7:0] _T_768 = _T_53 ? 8'h1 : _T_767; // @[Lookup.scala 33:37]
  wire [7:0] _T_769 = _T_51 ? 8'h1 : _T_768; // @[Lookup.scala 33:37]
  wire [7:0] _T_770 = _T_49 ? 8'h1 : _T_769; // @[Lookup.scala 33:37]
  wire [7:0] _T_771 = _T_47 ? 8'h1 : _T_770; // @[Lookup.scala 33:37]
  wire [7:0] _T_772 = _T_45 ? 8'h1 : _T_771; // @[Lookup.scala 33:37]
  wire [7:0] _T_773 = _T_43 ? 8'h1 : _T_772; // @[Lookup.scala 33:37]
  wire [7:0] _T_774 = _T_41 ? 8'h1 : _T_773; // @[Lookup.scala 33:37]
  wire [7:0] _T_775 = _T_39 ? 8'h1 : _T_774; // @[Lookup.scala 33:37]
  wire [7:0] _T_776 = _T_37 ? 8'h1 : _T_775; // @[Lookup.scala 33:37]
  wire [7:0] _T_777 = _T_35 ? 8'h1 : _T_776; // @[Lookup.scala 33:37]
  wire [7:0] _T_778 = _T_33 ? 8'h1 : _T_777; // @[Lookup.scala 33:37]
  wire [7:0] _T_779 = _T_31 ? 8'h1 : _T_778; // @[Lookup.scala 33:37]
  wire [7:0] _T_780 = _T_29 ? 8'h1 : _T_779; // @[Lookup.scala 33:37]
  wire [7:0] _T_781 = _T_25 ? 8'h1 : _T_780; // @[Lookup.scala 33:37]
  wire [7:0] _T_782 = _T_25 ? 8'h1 : _T_781; // @[Lookup.scala 33:37]
  wire [7:0] _T_783 = _T_23 ? 8'h1 : _T_782; // @[Lookup.scala 33:37]
  wire [7:0] _T_784 = _T_21 ? 8'h1 : _T_783; // @[Lookup.scala 33:37]
  wire [7:0] _T_785 = _T_19 ? 8'h1 : _T_784; // @[Lookup.scala 33:37]
  wire [7:0] _T_786 = _T_17 ? 8'h1 : _T_785; // @[Lookup.scala 33:37]
  wire [7:0] _T_787 = _T_15 ? 8'h1 : _T_786; // @[Lookup.scala 33:37]
  wire [7:0] _T_788 = _T_13 ? 8'h1 : _T_787; // @[Lookup.scala 33:37]
  wire [7:0] _T_789 = _T_11 ? 8'h1 : _T_788; // @[Lookup.scala 33:37]
  wire [7:0] _T_790 = _T_9 ? 8'h1 : _T_789; // @[Lookup.scala 33:37]
  wire [7:0] _T_791 = _T_7 ? 8'h1 : _T_790; // @[Lookup.scala 33:37]
  wire [7:0] _T_792 = _T_5 ? 8'h1 : _T_791; // @[Lookup.scala 33:37]
  wire [7:0] _T_793 = _T_3 ? 8'h1 : _T_792; // @[Lookup.scala 33:37]
  wire  _T_858 = _T_17 ? 1'h0 : _T_641; // @[Lookup.scala 33:37]
  wire  _T_859 = _T_15 ? 1'h0 : _T_858; // @[Lookup.scala 33:37]
  wire  _T_860 = _T_13 ? 1'h0 : _T_859; // @[Lookup.scala 33:37]
  wire  _T_861 = _T_11 ? 1'h0 : _T_860; // @[Lookup.scala 33:37]
  wire  _T_862 = _T_9 ? 1'h0 : _T_861; // @[Lookup.scala 33:37]
  wire  _T_863 = _T_7 ? 1'h0 : _T_862; // @[Lookup.scala 33:37]
  wire  _T_864 = _T_5 ? 1'h0 : _T_863; // @[Lookup.scala 33:37]
  wire  _T_865 = _T_3 ? 1'h0 : _T_864; // @[Lookup.scala 33:37]
  wire [1:0] _T_886 = _T_105 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_887 = _T_103 ? 2'h3 : _T_886; // @[Lookup.scala 33:37]
  wire [1:0] _T_888 = _T_101 ? 2'h3 : _T_887; // @[Lookup.scala 33:37]
  wire [1:0] _T_889 = _T_99 ? 2'h3 : _T_888; // @[Lookup.scala 33:37]
  wire [1:0] _T_890 = _T_97 ? 2'h3 : _T_889; // @[Lookup.scala 33:37]
  wire [1:0] _T_891 = _T_95 ? 2'h3 : _T_890; // @[Lookup.scala 33:37]
  wire [1:0] _T_892 = _T_93 ? 2'h0 : _T_891; // @[Lookup.scala 33:37]
  wire [1:0] _T_893 = _T_91 ? 2'h0 : _T_892; // @[Lookup.scala 33:37]
  wire [1:0] _T_894 = _T_89 ? 2'h0 : _T_893; // @[Lookup.scala 33:37]
  wire [1:0] _T_895 = _T_87 ? 2'h0 : _T_894; // @[Lookup.scala 33:37]
  wire [1:0] _T_896 = _T_85 ? 2'h0 : _T_895; // @[Lookup.scala 33:37]
  wire [1:0] _T_897 = _T_83 ? 2'h0 : _T_896; // @[Lookup.scala 33:37]
  wire [1:0] _T_898 = _T_81 ? 2'h0 : _T_897; // @[Lookup.scala 33:37]
  wire [1:0] _T_899 = _T_79 ? 2'h0 : _T_898; // @[Lookup.scala 33:37]
  wire [1:0] _T_900 = _T_77 ? 2'h0 : _T_899; // @[Lookup.scala 33:37]
  wire [1:0] _T_901 = _T_75 ? 2'h0 : _T_900; // @[Lookup.scala 33:37]
  wire [1:0] _T_902 = _T_73 ? 2'h0 : _T_901; // @[Lookup.scala 33:37]
  wire [1:0] _T_903 = _T_71 ? 2'h0 : _T_902; // @[Lookup.scala 33:37]
  wire [1:0] _T_904 = _T_69 ? 2'h0 : _T_903; // @[Lookup.scala 33:37]
  wire [1:0] _T_905 = _T_67 ? 2'h0 : _T_904; // @[Lookup.scala 33:37]
  wire [1:0] _T_906 = _T_65 ? 2'h0 : _T_905; // @[Lookup.scala 33:37]
  wire [1:0] _T_907 = _T_63 ? 2'h0 : _T_906; // @[Lookup.scala 33:37]
  wire [1:0] _T_908 = _T_61 ? 2'h0 : _T_907; // @[Lookup.scala 33:37]
  wire [1:0] _T_909 = _T_59 ? 2'h0 : _T_908; // @[Lookup.scala 33:37]
  wire [1:0] _T_910 = _T_57 ? 2'h0 : _T_909; // @[Lookup.scala 33:37]
  wire [1:0] _T_911 = _T_55 ? 2'h0 : _T_910; // @[Lookup.scala 33:37]
  wire [1:0] _T_912 = _T_53 ? 2'h0 : _T_911; // @[Lookup.scala 33:37]
  wire [1:0] _T_913 = _T_51 ? 2'h0 : _T_912; // @[Lookup.scala 33:37]
  wire [1:0] _T_914 = _T_49 ? 2'h0 : _T_913; // @[Lookup.scala 33:37]
  wire [1:0] _T_915 = _T_47 ? 2'h0 : _T_914; // @[Lookup.scala 33:37]
  wire [1:0] _T_916 = _T_45 ? 2'h0 : _T_915; // @[Lookup.scala 33:37]
  wire [1:0] _T_917 = _T_43 ? 2'h0 : _T_916; // @[Lookup.scala 33:37]
  wire [1:0] _T_918 = _T_41 ? 2'h0 : _T_917; // @[Lookup.scala 33:37]
  wire [1:0] _T_919 = _T_39 ? 2'h0 : _T_918; // @[Lookup.scala 33:37]
  wire [1:0] _T_920 = _T_37 ? 2'h0 : _T_919; // @[Lookup.scala 33:37]
  wire [1:0] _T_921 = _T_35 ? 2'h0 : _T_920; // @[Lookup.scala 33:37]
  wire [1:0] _T_922 = _T_33 ? 2'h0 : _T_921; // @[Lookup.scala 33:37]
  wire [1:0] _T_923 = _T_31 ? 2'h0 : _T_922; // @[Lookup.scala 33:37]
  wire [1:0] _T_924 = _T_29 ? 2'h0 : _T_923; // @[Lookup.scala 33:37]
  wire [1:0] _T_925 = _T_25 ? 2'h0 : _T_924; // @[Lookup.scala 33:37]
  wire [1:0] _T_926 = _T_25 ? 2'h0 : _T_925; // @[Lookup.scala 33:37]
  wire [1:0] _T_927 = _T_23 ? 2'h0 : _T_926; // @[Lookup.scala 33:37]
  wire [1:0] _T_928 = _T_21 ? 2'h0 : _T_927; // @[Lookup.scala 33:37]
  wire [1:0] _T_929 = _T_19 ? 2'h0 : _T_928; // @[Lookup.scala 33:37]
  wire [1:0] _T_930 = _T_17 ? 2'h1 : _T_929; // @[Lookup.scala 33:37]
  wire [1:0] _T_931 = _T_15 ? 2'h1 : _T_930; // @[Lookup.scala 33:37]
  wire [1:0] _T_932 = _T_13 ? 2'h1 : _T_931; // @[Lookup.scala 33:37]
  wire [1:0] _T_933 = _T_11 ? 2'h1 : _T_932; // @[Lookup.scala 33:37]
  wire [1:0] _T_934 = _T_9 ? 2'h1 : _T_933; // @[Lookup.scala 33:37]
  wire [1:0] _T_935 = _T_7 ? 2'h1 : _T_934; // @[Lookup.scala 33:37]
  wire [1:0] _T_936 = _T_5 ? 2'h1 : _T_935; // @[Lookup.scala 33:37]
  wire [1:0] _T_937 = _T_3 ? 2'h2 : _T_936; // @[Lookup.scala 33:37]
  wire [2:0] _T_953 = _T_115 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_954 = _T_113 ? 3'h5 : _T_953; // @[Lookup.scala 33:37]
  wire [2:0] _T_955 = _T_111 ? 3'h0 : _T_954; // @[Lookup.scala 33:37]
  wire [2:0] _T_956 = _T_109 ? 3'h5 : _T_955; // @[Lookup.scala 33:37]
  wire [2:0] _T_957 = _T_107 ? 3'h5 : _T_956; // @[Lookup.scala 33:37]
  wire [2:0] _T_958 = _T_105 ? 3'h2 : _T_957; // @[Lookup.scala 33:37]
  wire [2:0] _T_959 = _T_103 ? 3'h2 : _T_958; // @[Lookup.scala 33:37]
  wire [2:0] _T_960 = _T_101 ? 3'h4 : _T_959; // @[Lookup.scala 33:37]
  wire [2:0] _T_961 = _T_99 ? 3'h4 : _T_960; // @[Lookup.scala 33:37]
  wire [2:0] _T_962 = _T_97 ? 3'h3 : _T_961; // @[Lookup.scala 33:37]
  wire [2:0] _T_963 = _T_95 ? 3'h3 : _T_962; // @[Lookup.scala 33:37]
  wire [2:0] _T_964 = _T_93 ? 3'h0 : _T_963; // @[Lookup.scala 33:37]
  wire [2:0] _T_965 = _T_91 ? 3'h0 : _T_964; // @[Lookup.scala 33:37]
  wire [2:0] _T_966 = _T_89 ? 3'h0 : _T_965; // @[Lookup.scala 33:37]
  wire [2:0] _T_967 = _T_87 ? 3'h0 : _T_966; // @[Lookup.scala 33:37]
  wire [2:0] _T_968 = _T_85 ? 3'h0 : _T_967; // @[Lookup.scala 33:37]
  wire [2:0] _T_969 = _T_83 ? 3'h0 : _T_968; // @[Lookup.scala 33:37]
  wire [2:0] _T_970 = _T_81 ? 3'h0 : _T_969; // @[Lookup.scala 33:37]
  wire [2:0] _T_971 = _T_79 ? 3'h0 : _T_970; // @[Lookup.scala 33:37]
  wire [2:0] _T_972 = _T_77 ? 3'h0 : _T_971; // @[Lookup.scala 33:37]
  wire [2:0] _T_973 = _T_75 ? 3'h0 : _T_972; // @[Lookup.scala 33:37]
  wire [2:0] _T_974 = _T_73 ? 3'h0 : _T_973; // @[Lookup.scala 33:37]
  wire [2:0] _T_975 = _T_71 ? 3'h0 : _T_974; // @[Lookup.scala 33:37]
  wire [2:0] _T_976 = _T_69 ? 3'h0 : _T_975; // @[Lookup.scala 33:37]
  wire [2:0] _T_977 = _T_67 ? 3'h0 : _T_976; // @[Lookup.scala 33:37]
  wire [2:0] _T_978 = _T_65 ? 3'h0 : _T_977; // @[Lookup.scala 33:37]
  wire [2:0] _T_979 = _T_63 ? 3'h0 : _T_978; // @[Lookup.scala 33:37]
  wire [2:0] _T_980 = _T_61 ? 3'h0 : _T_979; // @[Lookup.scala 33:37]
  wire [2:0] _T_981 = _T_59 ? 3'h0 : _T_980; // @[Lookup.scala 33:37]
  wire [2:0] _T_982 = _T_57 ? 3'h0 : _T_981; // @[Lookup.scala 33:37]
  wire [2:0] _T_983 = _T_55 ? 3'h0 : _T_982; // @[Lookup.scala 33:37]
  wire [2:0] _T_984 = _T_53 ? 3'h0 : _T_983; // @[Lookup.scala 33:37]
  wire [2:0] _T_985 = _T_51 ? 3'h0 : _T_984; // @[Lookup.scala 33:37]
  wire [2:0] _T_986 = _T_49 ? 3'h0 : _T_985; // @[Lookup.scala 33:37]
  wire [2:0] _T_987 = _T_47 ? 3'h0 : _T_986; // @[Lookup.scala 33:37]
  wire [2:0] _T_988 = _T_45 ? 3'h0 : _T_987; // @[Lookup.scala 33:37]
  wire [2:0] _T_989 = _T_43 ? 3'h0 : _T_988; // @[Lookup.scala 33:37]
  wire [2:0] _T_990 = _T_41 ? 3'h0 : _T_989; // @[Lookup.scala 33:37]
  wire [2:0] _T_991 = _T_39 ? 3'h0 : _T_990; // @[Lookup.scala 33:37]
  wire [2:0] _T_992 = _T_37 ? 3'h0 : _T_991; // @[Lookup.scala 33:37]
  wire [2:0] _T_993 = _T_35 ? 3'h0 : _T_992; // @[Lookup.scala 33:37]
  wire [2:0] _T_994 = _T_33 ? 3'h0 : _T_993; // @[Lookup.scala 33:37]
  wire [2:0] _T_995 = _T_31 ? 3'h0 : _T_994; // @[Lookup.scala 33:37]
  wire [2:0] _T_996 = _T_29 ? 3'h0 : _T_995; // @[Lookup.scala 33:37]
  wire [2:0] _T_997 = _T_25 ? 3'h0 : _T_996; // @[Lookup.scala 33:37]
  wire [2:0] _T_998 = _T_25 ? 3'h0 : _T_997; // @[Lookup.scala 33:37]
  wire [2:0] _T_999 = _T_23 ? 3'h0 : _T_998; // @[Lookup.scala 33:37]
  wire [2:0] _T_1000 = _T_21 ? 3'h0 : _T_999; // @[Lookup.scala 33:37]
  wire [2:0] _T_1001 = _T_19 ? 3'h0 : _T_1000; // @[Lookup.scala 33:37]
  wire [2:0] _T_1002 = _T_17 ? 3'h0 : _T_1001; // @[Lookup.scala 33:37]
  wire [2:0] _T_1003 = _T_15 ? 3'h0 : _T_1002; // @[Lookup.scala 33:37]
  wire [2:0] _T_1004 = _T_13 ? 3'h0 : _T_1003; // @[Lookup.scala 33:37]
  wire [2:0] _T_1005 = _T_11 ? 3'h0 : _T_1004; // @[Lookup.scala 33:37]
  wire [2:0] _T_1006 = _T_9 ? 3'h0 : _T_1005; // @[Lookup.scala 33:37]
  wire [2:0] _T_1007 = _T_7 ? 3'h0 : _T_1006; // @[Lookup.scala 33:37]
  wire [2:0] _T_1008 = _T_5 ? 3'h0 : _T_1007; // @[Lookup.scala 33:37]
  wire [2:0] _T_1009 = _T_3 ? 3'h0 : _T_1008; // @[Lookup.scala 33:37]
  wire [2:0] _T_1010 = _T_145 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_1011 = _T_143 ? 3'h5 : _T_1010; // @[Lookup.scala 33:37]
  wire [2:0] _T_1012 = _T_141 ? 3'h0 : _T_1011; // @[Lookup.scala 33:37]
  wire [2:0] _T_1013 = _T_139 ? 3'h0 : _T_1012; // @[Lookup.scala 33:37]
  wire [2:0] _T_1014 = _T_137 ? 3'h5 : _T_1013; // @[Lookup.scala 33:37]
  wire [2:0] _T_1015 = _T_135 ? 3'h5 : _T_1014; // @[Lookup.scala 33:37]
  wire [2:0] _T_1016 = _T_133 ? 3'h0 : _T_1015; // @[Lookup.scala 33:37]
  wire [2:0] _T_1017 = _T_131 ? 3'h0 : _T_1016; // @[Lookup.scala 33:37]
  wire [2:0] _T_1018 = _T_129 ? 3'h5 : _T_1017; // @[Lookup.scala 33:37]
  wire [2:0] _T_1019 = _T_127 ? 3'h0 : _T_1018; // @[Lookup.scala 33:37]
  wire [2:0] _T_1020 = _T_125 ? 3'h0 : _T_1019; // @[Lookup.scala 33:37]
  wire [2:0] _T_1021 = _T_123 ? 3'h0 : _T_1020; // @[Lookup.scala 33:37]
  wire [2:0] _T_1022 = _T_121 ? 3'h0 : _T_1021; // @[Lookup.scala 33:37]
  wire [2:0] _T_1023 = _T_119 ? 3'h0 : _T_1022; // @[Lookup.scala 33:37]
  wire [2:0] _T_1024 = _T_117 ? 3'h0 : _T_1023; // @[Lookup.scala 33:37]
  wire [2:0] _T_1025 = _T_115 ? 3'h0 : _T_1024; // @[Lookup.scala 33:37]
  wire [2:0] _T_1026 = _T_113 ? 3'h0 : _T_1025; // @[Lookup.scala 33:37]
  wire [2:0] _T_1027 = _T_111 ? 3'h0 : _T_1026; // @[Lookup.scala 33:37]
  wire [2:0] _T_1028 = _T_109 ? 3'h0 : _T_1027; // @[Lookup.scala 33:37]
  wire [2:0] _T_1029 = _T_107 ? 3'h0 : _T_1028; // @[Lookup.scala 33:37]
  wire [2:0] _T_1030 = _T_105 ? 3'h0 : _T_1029; // @[Lookup.scala 33:37]
  wire [2:0] _T_1031 = _T_103 ? 3'h0 : _T_1030; // @[Lookup.scala 33:37]
  wire [2:0] _T_1032 = _T_101 ? 3'h0 : _T_1031; // @[Lookup.scala 33:37]
  wire [2:0] _T_1033 = _T_99 ? 3'h0 : _T_1032; // @[Lookup.scala 33:37]
  wire [2:0] _T_1034 = _T_97 ? 3'h0 : _T_1033; // @[Lookup.scala 33:37]
  wire [2:0] _T_1035 = _T_95 ? 3'h0 : _T_1034; // @[Lookup.scala 33:37]
  wire [2:0] _T_1036 = _T_93 ? 3'h0 : _T_1035; // @[Lookup.scala 33:37]
  wire [2:0] _T_1037 = _T_91 ? 3'h0 : _T_1036; // @[Lookup.scala 33:37]
  wire [2:0] _T_1038 = _T_89 ? 3'h0 : _T_1037; // @[Lookup.scala 33:37]
  wire [2:0] _T_1039 = _T_87 ? 3'h0 : _T_1038; // @[Lookup.scala 33:37]
  wire [2:0] _T_1040 = _T_85 ? 3'h0 : _T_1039; // @[Lookup.scala 33:37]
  wire [2:0] _T_1041 = _T_83 ? 3'h0 : _T_1040; // @[Lookup.scala 33:37]
  wire [2:0] _T_1042 = _T_81 ? 3'h0 : _T_1041; // @[Lookup.scala 33:37]
  wire [2:0] _T_1043 = _T_79 ? 3'h0 : _T_1042; // @[Lookup.scala 33:37]
  wire [2:0] _T_1044 = _T_77 ? 3'h0 : _T_1043; // @[Lookup.scala 33:37]
  wire [2:0] _T_1045 = _T_75 ? 3'h0 : _T_1044; // @[Lookup.scala 33:37]
  wire [2:0] _T_1046 = _T_73 ? 3'h0 : _T_1045; // @[Lookup.scala 33:37]
  wire [2:0] _T_1047 = _T_71 ? 3'h0 : _T_1046; // @[Lookup.scala 33:37]
  wire [2:0] _T_1048 = _T_69 ? 3'h5 : _T_1047; // @[Lookup.scala 33:37]
  wire [2:0] _T_1049 = _T_67 ? 3'h5 : _T_1048; // @[Lookup.scala 33:37]
  wire [2:0] _T_1050 = _T_65 ? 3'h0 : _T_1049; // @[Lookup.scala 33:37]
  wire [2:0] _T_1051 = _T_63 ? 3'h0 : _T_1050; // @[Lookup.scala 33:37]
  wire [2:0] _T_1052 = _T_61 ? 3'h0 : _T_1051; // @[Lookup.scala 33:37]
  wire [2:0] _T_1053 = _T_59 ? 3'h0 : _T_1052; // @[Lookup.scala 33:37]
  wire [2:0] _T_1054 = _T_57 ? 3'h5 : _T_1053; // @[Lookup.scala 33:37]
  wire [2:0] _T_1055 = _T_55 ? 3'h0 : _T_1054; // @[Lookup.scala 33:37]
  wire [2:0] _T_1056 = _T_53 ? 3'h5 : _T_1055; // @[Lookup.scala 33:37]
  wire [2:0] _T_1057 = _T_51 ? 3'h5 : _T_1056; // @[Lookup.scala 33:37]
  wire [2:0] _T_1058 = _T_49 ? 3'h0 : _T_1057; // @[Lookup.scala 33:37]
  wire [2:0] _T_1059 = _T_47 ? 3'h0 : _T_1058; // @[Lookup.scala 33:37]
  wire [2:0] _T_1060 = _T_45 ? 3'h5 : _T_1059; // @[Lookup.scala 33:37]
  wire [2:0] _T_1061 = _T_43 ? 3'h5 : _T_1060; // @[Lookup.scala 33:37]
  wire [2:0] _T_1062 = _T_41 ? 3'h0 : _T_1061; // @[Lookup.scala 33:37]
  wire [2:0] _T_1063 = _T_39 ? 3'h0 : _T_1062; // @[Lookup.scala 33:37]
  wire [2:0] _T_1064 = _T_37 ? 3'h0 : _T_1063; // @[Lookup.scala 33:37]
  wire [2:0] _T_1065 = _T_35 ? 3'h0 : _T_1064; // @[Lookup.scala 33:37]
  wire [2:0] _T_1066 = _T_33 ? 3'h0 : _T_1065; // @[Lookup.scala 33:37]
  wire [2:0] _T_1067 = _T_31 ? 3'h0 : _T_1066; // @[Lookup.scala 33:37]
  wire [2:0] _T_1068 = _T_29 ? 3'h5 : _T_1067; // @[Lookup.scala 33:37]
  wire [2:0] _T_1069 = _T_25 ? 3'h5 : _T_1068; // @[Lookup.scala 33:37]
  wire [2:0] _T_1070 = _T_25 ? 3'h0 : _T_1069; // @[Lookup.scala 33:37]
  wire [2:0] _T_1071 = _T_23 ? 3'h0 : _T_1070; // @[Lookup.scala 33:37]
  wire [2:0] _T_1072 = _T_21 ? 3'h0 : _T_1071; // @[Lookup.scala 33:37]
  wire [2:0] _T_1073 = _T_19 ? 3'h0 : _T_1072; // @[Lookup.scala 33:37]
  wire [2:0] _T_1074 = _T_17 ? 3'h0 : _T_1073; // @[Lookup.scala 33:37]
  wire [2:0] _T_1075 = _T_15 ? 3'h0 : _T_1074; // @[Lookup.scala 33:37]
  wire [2:0] _T_1076 = _T_13 ? 3'h0 : _T_1075; // @[Lookup.scala 33:37]
  wire [2:0] _T_1077 = _T_11 ? 3'h0 : _T_1076; // @[Lookup.scala 33:37]
  wire [2:0] _T_1078 = _T_9 ? 3'h0 : _T_1077; // @[Lookup.scala 33:37]
  wire [2:0] _T_1079 = _T_7 ? 3'h0 : _T_1078; // @[Lookup.scala 33:37]
  wire [2:0] _T_1080 = _T_5 ? 3'h0 : _T_1079; // @[Lookup.scala 33:37]
  wire [2:0] _T_1081 = _T_3 ? 3'h0 : _T_1080; // @[Lookup.scala 33:37]
  wire  _T_1117 = ~cs_valid_inst; // @[cpath.scala 163:46]
  wire  temp_exception = io_imem_resp_valid & _T_1117; // @[cpath.scala 163:43]
  wire  _T_1082 = temp_exception | io_d2c_isredir; // @[cpath.scala 146:25]
  wire  _T_1083 = cs_branch == 4'h0; // @[cpath.scala 147:20]
  wire  _T_1084 = cs_branch == 4'h1; // @[cpath.scala 148:20]
  wire [2:0] _T_1085 = io_d2c_iseq ? 3'h2 : 3'h0; // @[cpath.scala 148:38]
  wire  _T_1086 = cs_branch == 4'h2; // @[cpath.scala 149:20]
  wire  _T_1087 = ~io_d2c_iseq; // @[cpath.scala 149:40]
  wire [2:0] _T_1088 = _T_1087 ? 3'h2 : 3'h0; // @[cpath.scala 149:39]
  wire  _T_1089 = cs_branch == 4'h5; // @[cpath.scala 150:20]
  wire  _T_1090 = ~io_d2c_islt; // @[cpath.scala 150:39]
  wire [2:0] _T_1091 = _T_1090 ? 3'h2 : 3'h0; // @[cpath.scala 150:38]
  wire  _T_1092 = cs_branch == 4'h6; // @[cpath.scala 151:20]
  wire  _T_1093 = ~io_d2c_isltu; // @[cpath.scala 151:40]
  wire [2:0] _T_1094 = _T_1093 ? 3'h2 : 3'h0; // @[cpath.scala 151:39]
  wire  _T_1095 = cs_branch == 4'h3; // @[cpath.scala 152:20]
  wire [2:0] _T_1096 = io_d2c_islt ? 3'h2 : 3'h0; // @[cpath.scala 152:38]
  wire  _T_1097 = cs_branch == 4'h4; // @[cpath.scala 153:20]
  wire [2:0] _T_1098 = io_d2c_isltu ? 3'h2 : 3'h0; // @[cpath.scala 153:39]
  wire  _T_1099 = cs_branch == 4'h7; // @[cpath.scala 154:20]
  wire  _T_1100 = cs_branch == 4'h8; // @[cpath.scala 155:20]
  wire [2:0] _T_1101 = _T_1100 ? 3'h3 : 3'h0; // @[Mux.scala 98:16]
  wire [2:0] _T_1102 = _T_1099 ? 3'h1 : _T_1101; // @[Mux.scala 98:16]
  wire [2:0] _T_1103 = _T_1097 ? _T_1098 : _T_1102; // @[Mux.scala 98:16]
  wire [2:0] _T_1104 = _T_1095 ? _T_1096 : _T_1103; // @[Mux.scala 98:16]
  wire [2:0] _T_1105 = _T_1092 ? _T_1094 : _T_1104; // @[Mux.scala 98:16]
  wire [2:0] _T_1106 = _T_1089 ? _T_1091 : _T_1105; // @[Mux.scala 98:16]
  wire [2:0] _T_1107 = _T_1086 ? _T_1088 : _T_1106; // @[Mux.scala 98:16]
  wire [2:0] _T_1108 = _T_1084 ? _T_1085 : _T_1107; // @[Mux.scala 98:16]
  wire [2:0] _T_1109 = _T_1083 ? 3'h0 : _T_1108; // @[Mux.scala 98:16]
  wire [2:0] _T_1110 = _T_1082 ? 3'h4 : _T_1109; // @[Mux.scala 98:16]
  wire [1:0] temp_pc_sel = _T_1110[1:0]; // @[cpath.scala 141:27 cpath.scala 145:17]
  assign io_c2d_cp_pc_sel = {{1'd0}, temp_pc_sel}; // @[cpath.scala 179:33]
  assign io_c2d_cp_op1_sel = _T_1 ? 2'h0 : _T_361; // @[cpath.scala 180:33]
  assign io_c2d_cp_op2_sel = _T_1 ? 2'h0 : _T_433; // @[cpath.scala 181:33]
  assign io_c2d_cp_alu_sel = _T_1 ? 5'h0 : _T_505; // @[cpath.scala 182:33]
  assign io_c2d_cp_reg_wen = _T_1 ? 1'h0 : _T_577; // @[cpath.scala 183:33]
  assign io_c2d_cp_mem_en = _T_1 ? 1'h0 : _T_649; // @[cpath.scala 184:33]
  assign io_c2d_cp_mem_read_op = _T_1 ? 3'h0 : _T_721; // @[cpath.scala 185:33]
  assign io_c2d_cp_mem_write_mask = _T_1 ? 8'h1 : _T_793; // @[cpath.scala 186:33]
  assign io_c2d_cp_mem_wen = _T_1 ? 1'h0 : _T_865; // @[cpath.scala 187:33]
  assign io_c2d_cp_alu_ext_sel = _T_1 ? 3'h0 : _T_1081; // @[cpath.scala 188:33]
  assign io_c2d_cp_wb_sel = _T_1 ? 2'h2 : _T_937; // @[cpath.scala 189:33]
  assign io_c2d_cp_csr_op = _T_1 ? 3'h0 : _T_1009; // @[cpath.scala 190:33]
  assign io_c2d_hasexception = 1'h0;
  assign io_c2d_shouldstall = 1'h0;
  assign io_imem_req_ready = 1'h0;
  assign io_imem_resp_valid = 1'h0;
  assign io_imem_resp_bits_rdata = 64'h0;
  assign io_dmem_req_ready = 1'h0;
  assign io_dmem_resp_valid = 1'h0;
  assign io_dmem_resp_bits_rdata = 64'h0;
endmodule
