module alu_module(
  input         clock,
  input         reset,
  input  [63:0] io_input1,
  input  [63:0] io_input2,
  input  [4:0]  io_op,
  input  [2:0]  io_res_ext_op,
  output [63:0] io_res
);
  wire [63:0] add_res = io_input1 + io_input2; // @[alu.scala 29:26]
  wire [5:0] sham = io_input2[5:0]; // @[alu.scala 31:25]
  wire  _T_2 = io_op == 5'h0; // @[alu.scala 36:16]
  wire  _T_3 = io_op == 5'h1; // @[alu.scala 37:16]
  wire [63:0] _T_5 = io_input1 - io_input2; // @[alu.scala 37:43]
  wire  _T_6 = io_op == 5'h2; // @[alu.scala 38:16]
  wire [63:0] _T_7 = io_input1 & io_input2; // @[alu.scala 38:43]
  wire  _T_8 = io_op == 5'h3; // @[alu.scala 39:16]
  wire [63:0] _T_9 = io_input1 | io_input2; // @[alu.scala 39:42]
  wire  _T_10 = io_op == 5'h4; // @[alu.scala 40:16]
  wire [63:0] _T_11 = io_input1 ^ io_input2; // @[alu.scala 40:43]
  wire  _T_12 = io_op == 5'h5; // @[alu.scala 41:16]
  wire [126:0] _GEN_0 = {{63'd0}, io_input1}; // @[alu.scala 41:44]
  wire [126:0] _T_13 = _GEN_0 << sham; // @[alu.scala 41:44]
  wire  _T_15 = io_op == 5'h6; // @[alu.scala 42:16]
  wire [63:0] _T_16 = io_input1; // @[alu.scala 42:49]
  wire  _T_18 = $signed(io_input1) < $signed(io_input2); // @[alu.scala 42:52]
  wire  _T_19 = io_op == 5'h7; // @[alu.scala 43:16]
  wire  _T_20 = io_input1 < io_input2; // @[alu.scala 43:53]
  wire  _T_21 = io_op == 5'h8; // @[alu.scala 44:16]
  wire [63:0] _T_24 = $signed(io_input1) >>> sham; // @[alu.scala 44:68]
  wire  _T_25 = io_op == 5'h9; // @[alu.scala 45:16]
  wire [31:0] _T_27 = io_input1[31:0]; // @[alu.scala 45:57]
  wire [31:0] _T_29 = $signed(_T_27) >>> sham; // @[alu.scala 45:75]
  wire  _T_30 = io_op == 5'ha; // @[alu.scala 46:16]
  wire [63:0] _T_31 = io_input1 >> sham; // @[alu.scala 46:53]
  wire  _T_32 = io_op == 5'hb; // @[alu.scala 47:16]
  wire [31:0] _T_34 = io_input1[31:0] >> sham; // @[alu.scala 47:60]
  wire  _T_35 = io_op == 5'hc; // @[alu.scala 48:16]
  wire  _T_36 = io_op == 5'hd; // @[alu.scala 49:16]
  wire [127:0] _T_39 = $signed(io_input1) * $signed(io_input2); // @[alu.scala 49:53]
  wire  _T_41 = io_op == 5'he; // @[alu.scala 50:16]
  wire  _T_46 = io_op == 5'hf; // @[alu.scala 51:16]
  wire [64:0] _T_49 = {1'h0,io_input2}; // @[alu.scala 51:88]
  wire [64:0] _GEN_1 = {{1{_T_16[63]}},_T_16}; // @[alu.scala 51:56]
  wire [128:0] _T_50 = $signed(_GEN_1) * $signed(_T_49); // @[alu.scala 51:56]
  wire  _T_52 = io_op == 5'h10; // @[alu.scala 52:16]
  wire [127:0] _T_53 = io_input1 * io_input2; // @[alu.scala 52:55]
  wire  _T_55 = io_op == 5'h11; // @[alu.scala 53:16]
  wire [63:0] _T_59 = $signed(io_input1) % $signed(io_input2); // @[alu.scala 53:81]
  wire  _T_60 = io_op == 5'h12; // @[alu.scala 54:16]
  wire [63:0] _GEN_2 = io_input1 % io_input2; // @[alu.scala 54:54]
  wire [63:0] _T_61 = _GEN_2[63:0]; // @[alu.scala 54:54]
  wire  _T_62 = io_op == 5'h13; // @[alu.scala 55:16]
  wire [31:0] _GEN_3 = io_input1[31:0] % io_input2[31:0]; // @[alu.scala 55:61]
  wire [31:0] _T_65 = _GEN_3[31:0]; // @[alu.scala 55:61]
  wire  _T_66 = io_op == 5'h14; // @[alu.scala 56:16]
  wire [31:0] _T_70 = io_input2[31:0]; // @[alu.scala 56:84]
  wire [31:0] _T_72 = $signed(_T_27) % $signed(_T_70); // @[alu.scala 56:94]
  wire  _T_73 = io_op == 5'h15; // @[alu.scala 57:16]
  wire [64:0] _T_77 = $signed(io_input1) / $signed(io_input2); // @[alu.scala 57:81]
  wire  _T_78 = io_op == 5'h16; // @[alu.scala 58:16]
  wire [31:0] _T_81 = io_input1[31:0] / io_input2[31:0]; // @[alu.scala 58:61]
  wire  _T_82 = io_op == 5'h17; // @[alu.scala 59:16]
  wire [32:0] _T_88 = $signed(_T_27) / $signed(_T_70); // @[alu.scala 59:94]
  wire [63:0] _T_89 = _T_82 ? {{31'd0}, _T_88} : add_res; // @[Mux.scala 98:16]
  wire [63:0] _T_90 = _T_78 ? {{32'd0}, _T_81} : _T_89; // @[Mux.scala 98:16]
  wire [64:0] _T_91 = _T_73 ? _T_77 : {{1'd0}, _T_90}; // @[Mux.scala 98:16]
  wire [64:0] _T_92 = _T_66 ? {{33'd0}, _T_72} : _T_91; // @[Mux.scala 98:16]
  wire [64:0] _T_93 = _T_62 ? {{33'd0}, _T_65} : _T_92; // @[Mux.scala 98:16]
  wire [64:0] _T_94 = _T_60 ? {{1'd0}, _T_61} : _T_93; // @[Mux.scala 98:16]
  wire [64:0] _T_95 = _T_55 ? {{1'd0}, _T_59} : _T_94; // @[Mux.scala 98:16]
  wire [64:0] _T_96 = _T_52 ? {{1'd0}, _T_53[127:64]} : _T_95; // @[Mux.scala 98:16]
  wire [64:0] _T_97 = _T_46 ? {{1'd0}, _T_50[127:64]} : _T_96; // @[Mux.scala 98:16]
  wire [64:0] _T_98 = _T_41 ? {{1'd0}, _T_39[127:64]} : _T_97; // @[Mux.scala 98:16]
  wire [64:0] _T_99 = _T_36 ? {{1'd0}, _T_39[63:0]} : _T_98; // @[Mux.scala 98:16]
  wire [64:0] _T_100 = _T_35 ? {{1'd0}, io_input1} : _T_99; // @[Mux.scala 98:16]
  wire [64:0] _T_101 = _T_32 ? {{33'd0}, _T_34} : _T_100; // @[Mux.scala 98:16]
  wire [64:0] _T_102 = _T_30 ? {{1'd0}, _T_31} : _T_101; // @[Mux.scala 98:16]
  wire [64:0] _T_103 = _T_25 ? {{33'd0}, _T_29} : _T_102; // @[Mux.scala 98:16]
  wire [64:0] _T_104 = _T_21 ? {{1'd0}, _T_24} : _T_103; // @[Mux.scala 98:16]
  wire [64:0] _T_105 = _T_19 ? {{64'd0}, _T_20} : _T_104; // @[Mux.scala 98:16]
  wire [64:0] _T_106 = _T_15 ? {{64'd0}, _T_18} : _T_105; // @[Mux.scala 98:16]
  wire [64:0] _T_107 = _T_12 ? {{1'd0}, _T_13[63:0]} : _T_106; // @[Mux.scala 98:16]
  wire [64:0] _T_108 = _T_10 ? {{1'd0}, _T_11} : _T_107; // @[Mux.scala 98:16]
  wire [64:0] _T_109 = _T_8 ? {{1'd0}, _T_9} : _T_108; // @[Mux.scala 98:16]
  wire [64:0] _T_110 = _T_6 ? {{1'd0}, _T_7} : _T_109; // @[Mux.scala 98:16]
  wire [64:0] _T_111 = _T_3 ? {{1'd0}, _T_5} : _T_110; // @[Mux.scala 98:16]
  wire [64:0] _T_112 = _T_2 ? {{1'd0}, add_res} : _T_111; // @[Mux.scala 98:16]
  wire  _T_113 = io_res_ext_op == 3'h0; // @[alu.scala 64:24]
  wire  _T_114 = io_res_ext_op == 3'h1; // @[alu.scala 65:24]
  wire [63:0] res_temp = _T_112[63:0]; // @[alu.scala 27:24 alu.scala 35:14]
  wire [55:0] _T_117 = res_temp[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_119 = {_T_117,res_temp[7:0]}; // @[Cat.scala 29:58]
  wire  _T_120 = io_res_ext_op == 3'h2; // @[alu.scala 66:24]
  wire [63:0] _T_123 = {56'h0,res_temp[7:0]}; // @[Cat.scala 29:58]
  wire  _T_124 = io_res_ext_op == 3'h3; // @[alu.scala 67:24]
  wire [47:0] _T_127 = res_temp[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_129 = {_T_127,res_temp[15:0]}; // @[Cat.scala 29:58]
  wire  _T_130 = io_res_ext_op == 3'h4; // @[alu.scala 68:24]
  wire [63:0] _T_133 = {48'h0,res_temp[15:0]}; // @[Cat.scala 29:58]
  wire  _T_134 = io_res_ext_op == 3'h5; // @[alu.scala 69:24]
  wire [31:0] _T_137 = res_temp[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_139 = {_T_137,res_temp[31:0]}; // @[Cat.scala 29:58]
  wire  _T_140 = io_res_ext_op == 3'h6; // @[alu.scala 70:24]
  wire [63:0] _T_143 = {32'h0,res_temp[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_144 = _T_140 ? _T_143 : res_temp; // @[Mux.scala 98:16]
  wire [63:0] _T_145 = _T_134 ? _T_139 : _T_144; // @[Mux.scala 98:16]
  wire [63:0] _T_146 = _T_130 ? _T_133 : _T_145; // @[Mux.scala 98:16]
  wire [63:0] _T_147 = _T_124 ? _T_129 : _T_146; // @[Mux.scala 98:16]
  wire [63:0] _T_148 = _T_120 ? _T_123 : _T_147; // @[Mux.scala 98:16]
  wire [63:0] _T_149 = _T_114 ? _T_119 : _T_148; // @[Mux.scala 98:16]
  assign io_res = _T_113 ? res_temp : _T_149; // @[alu.scala 63:12]
endmodule
